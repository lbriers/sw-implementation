--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"004124230031222300112023340111730000001300000013000000131140006f",
        INIT_01 => X"02c1242302b1222302a1202300912e2300812c2300712a230061282300512623",
        INIT_02 => X"05412423053122230521202303112e2303012c2302f12a2302e1282302d12623",
        INIT_03 => X"07c1242307b1222307a1202305912e2305812c2305712a230561282305512623",
        INIT_04 => X"00812203004121830001208371d000ef3420357307f12a2307e1282307d12623",
        INIT_05 => X"02812603024125830201250301c1248301812403014123830101230300c12283",
        INIT_06 => X"04812a03044129830401290303c1288303812803034127830301270302c12683",
        INIT_07 => X"06812e0306412d8306012d0305c12c8305812c0305412b8305012b0304c12a83",
        INIT_08 => X"000001930000011300000093302000733401117307412f8307012f0306c12e83",
        INIT_09 => X"0000059300000513000004930000041300000393000003130000029300000213",
        INIT_0A => X"0000099300000913000008930000081300000793000007130000069300000613",
        INIT_0B => X"00000d9300000d1300000c9300000c1300000b9300000b1300000a9300000a13",
        INIT_0C => X"0000113700018213eef18193deadc1b700000f9300000f1300000e9300000e13",
        INIT_0D => X"30411073fff001133004507330511073e6810113000001173401107300010113",
        INIT_0E => X"00112023ff4101130540006f605000ef0010007360d000effe01011300001137",
        INIT_0F => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_10 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_11 => X"0201041300812c2300112e23fe0101130000006f0000006f0000806700c10113",
        INIT_12 => X"fea42623679000effec4250300500593fef42623fe078793fec42783fea42623",
        INIT_13 => X"0181240301c1208300078513fec42783fea426236dd000effec4250300900593",
        INIT_14 => X"feb42423fea426230201041300812c2300112e23fe0101130000806702010113",
        INIT_15 => X"94e7aa23fe842703000047b794e7a823fec42703000047b7fed42023fec42223",
        INIT_16 => X"01c120830000001394e7ae23fe042703000047b794e7ac23fe442703000047b7",
        INIT_17 => X"000507930201041300812c2300112e23fe010113000080670201011301812403",
        INIT_18 => X"00f717b30037979340f687b3003006939607a783000047b7fef44703fef407a3",
        INIT_19 => X"9607a703000047b796e7a223000047b700f707339647a783000047b700078713",
        INIT_1A => X"9607a023000047b700e7a0239647270300004737800007b702f7146300300793",
        INIT_1B => X"96e7a023000047b7001787139607a783000047b701c0006f9607a223000047b7",
        INIT_1C => X"0281242302112623fd01011300008067020101130181240301c1208300000013",
        INIT_1D => X"000785130ff7f793fec42783fef426230187d793fdc42783fca42e2303010413",
        INIT_1E => X"000785130ff7f793fec42783fef426230ff7f7930107d793fdc42783f2dff0ef",
        INIT_1F => X"000785130ff7f793fec42783fef426230ff7f7930087d793fdc42783f0dff0ef",
        INIT_20 => X"ed1ff0ef000785130ff7f793fec42783fef426230ff7f793fdc42783eedff0ef",
        INIT_21 => X"0281242302112623fd01011300008067030101130281240302c1208300000013",
        INIT_22 => X"fef4262300f707b3fec4270301879793fdc42783fe042623fca42e2303010413",
        INIT_23 => X"fdc42783fef4262300f707b3fec4270300f777b300ff07b700879713fdc42783",
        INIT_24 => X"fdc42783fef4262300f707b3fec4270300f777b3f0078793000107b70087d713",
        INIT_25 => X"0281240302c1208300078513fec42783fef4262300f707b3fec427030187d793",
        INIT_26 => X"feb42423fea426230201041300812c2300112e23fe0101130000806703010113",
        INIT_27 => X"07100513d91ff0ef0000051300000593000006130ff00693fed42023fec42223",
        INIT_28 => X"fec42783148010ef06600513150010ef06900513158010ef06f00513160010ef",
        INIT_29 => X"000785130ff7f7930107d793fec42783134010ef000785130ff7f7930187d793",
        INIT_2A => X"0ff7f793fec4278310c010ef000785130ff7f7930087d793fec42783120010ef",
        INIT_2B => X"fe8427830e8010ef000785130ff7f7930187d793fe8427830fc010ef00078513",
        INIT_2C => X"000785130ff7f7930087d793fe8427830d4010ef000785130ff7f7930107d793",
        INIT_2D => X"000785130ff7f793fe4427830b0010ef000785130ff7f793fe8427830c0010ef",
        INIT_2E => X"0181240301c1208300000013090010ef000785130ff7f793fe0427830a0010ef",
        INIT_2F => X"feb42423fea42623030104130281242302112623fd0101130000806702010113",
        INIT_30 => X"fdc42783fec42703fd142823fd042a23fcf42c23fce42e23fed42023fec42223",
        INIT_31 => X"0300006f0000079300f70663fd842783fe8427030440006f0000079300f70663",
        INIT_32 => X"00f70663fd042783fe04270301c0006f0000079300f70663fd442783fe442703",
        INIT_33 => X"00008067030101130281240302c1208300078513001007930080006f00000793",
        INIT_34 => X"fcd42823fcc42a23fcb42c23fca42e23030104130281242302112623fd010113",
        INIT_35 => X"95c7a783000047b79587a603000047b79547a683000047b79507a703000047b7",
        INIT_36 => X"f0dff0effdc42503fd842583fd442603fd042683000687930006081300078893",
        INIT_37 => X"9687a783000047b704e7e86303f007939687a703000047b70607806300050793",
        INIT_38 => X"fd842703000047b794e7a823fdc42703000047b796e7a423000047b700178713",
        INIT_39 => X"0010079394e7ae23fd042703000047b794e7ac23fd442703000047b794e7aa23",
        INIT_3A => X"fef426230bf787939687a783000047b7020786639687a783000047b703c0006f",
        INIT_3B => X"00078513000007939607a423000047b76f5000ef000785130ff7f793fec42783",
        INIT_3C => X"00912a2300812c2300112e23fe01011300008067030101130281240302c12083",
        INIT_3D => X"a1dff0ef00300513fec42583fed42023fec42223feb42423fea4262302010413",
        INIT_3E => X"00700513fe44258300f484b300050793a0dff0ef00500513fe84258300050493",
        INIT_3F => X"00f487b3000507939e5ff0ef00b00513fe04258300f484b3000507939f9ff0ef",
        INIT_40 => X"fd0101130000806702010113014124830181240301c120830007851303f7f793",
        INIT_41 => X"fd042683fcd42823fcc42a23fcb42c23fca42e23030104130281242302112623",
        INIT_42 => X"fec4278355078713000037b7fea42623f45ff0effdc42503fd842583fd442603",
        INIT_43 => X"00f707b300479793fec4278355078713000037b70007a50300f707b300479793",
        INIT_44 => X"000037b70087a60300f707b300479793fec4278355078713000037b70047a583",
        INIT_45 => X"fd842783fd442803fd04288300c7a68300f707b300479793fec4278355078713",
        INIT_46 => X"fe842783fef4242303f7f793fec4278304078c6300050793d25ff0effdc42703",
        INIT_47 => X"fd842703000047b794e7a823fdc42703000047b7579000ef000785130ff7f793",
        INIT_48 => X"0010079394e7ae23fd042703000047b794e7ac23fd442703000047b794e7aa23",
        INIT_49 => X"00e7a023fdc4270300f707b300479793fec4278355078713000037b70780006f",
        INIT_4A => X"000037b700e7a223fd84270300f707b300479793fec4278355078713000037b7",
        INIT_4B => X"55078713000037b700e7a423fd44270300f707b300479793fec4278355078713",
        INIT_4C => X"02c12083000785130000079300e7a623fd04270300f707b300479793fec42783",
        INIT_4D => X"fca426230401041302812c2302112e23fc010113000080670301011302812403",
        INIT_4E => X"0027879340f707b3fcc427039507a783000047b7fcd42023fcc42223fcb42423",
        INIT_4F => X"0ff7f7930027879340f707b3fc8427039547a783000047b7fef426230ff7f793",
        INIT_50 => X"fef422230ff7f7930027879340f707b3fc4427039587a783000047b7fef42423",
        INIT_51 => X"00e7f66300300793fe8427030c40006f0000079300e7f66300300793fec42703",
        INIT_52 => X"fec4278309c0006f0000079300e7f66300300793fe4427030b00006f00000793",
        INIT_53 => X"fe442783fef4242300c7f79300279793fe842783fef426230307f79300479793",
        INIT_54 => X"fe44278300f70733fe842783fec42703fef4202304000793fef422230037f793",
        INIT_55 => X"3a5000ef000785130ff7f793fdc42783fcf42e2300f707b3fe04270300f707b3",
        INIT_56 => X"fc442703000047b794e7aa23fc842703000047b794e7a823fcc42703000047b7",
        INIT_57 => X"0381240303c12083000785130010079394e7ae23fc042703000047b794e7ac23",
        INIT_58 => X"fcb42c23fca42e23030104130281242302112623fd0101130000806704010113",
        INIT_59 => X"0ff7f7930207879340f707b3fd8427039547a783000047b7fcd42823fcc42a23",
        INIT_5A => X"9507a783000047b71180006f0000079300e7f66303f00793fec42703fef42623",
        INIT_5B => X"0087879300f707b340f687b3fd8427839547a683000047b740f70733fdc42703",
        INIT_5C => X"000047b70d40006f0000079300e7f66300f00793fe842703fef424230ff7f793",
        INIT_5D => X"00f707b340f687b3fd8427839547a683000047b740f70733fd4427039587a783",
        INIT_5E => X"0900006f0000079300e7f66300f00793fe442703fef422230ff7f79300878793",
        INIT_5F => X"fe042783fef4202300f707b3fe04270303f7f793fec42783fef4202308000793",
        INIT_60 => X"00f7f793fe4427830ff7f71300479793fe842783259000ef000785130ff7f793",
        INIT_61 => X"fdc42703000047b722d000ef000785130ff7f793fe042783fef4202300f707b3",
        INIT_62 => X"000047b794e7ac23fd442703000047b794e7aa23fd842703000047b794e7a823",
        INIT_63 => X"00008067030101130281240302c12083000785130010079394e7ae23fd042703",
        INIT_64 => X"fed42023fec42223feb42423fea426230201041300812c2300112e23fe010113",
        INIT_65 => X"0ff7f793fec427831ad000ef0fe0051306f71a63fe04270395c7a783000047b7",
        INIT_66 => X"0ff7f793fe44278318d000ef000785130ff7f793fe84278319d000ef00078513",
        INIT_67 => X"94e7aa23fe842703000047b794e7a823fec42703000047b717d000ef00078513",
        INIT_68 => X"0080006f0010079394e7ae23fe042703000047b794e7ac23fe442703000047b7",
        INIT_69 => X"00112e23fe01011300008067020101130181240301c120830007851300000793",
        INIT_6A => X"105000ef0ff00513fed42023fec42223feb42423fea426230201041300812c23",
        INIT_6B => X"0e5000ef000785130ff7f793fe8427830f5000ef000785130ff7f793fec42783",
        INIT_6C => X"0c5000ef000785130ff7f793fe0427830d5000ef000785130ff7f793fe442783",
        INIT_6D => X"00812c2300112e23fe01011300008067020101130181240301c1208300000013",
        INIT_6E => X"fff7879300f707b3fec427839687a703000047b7fef426230c00079302010413",
        INIT_6F => X"000005139607a423000047b7071000ef000785130ff7f793fe842783fef42423",
        INIT_70 => X"00000513049000ef00000513051000ef00000513059000ef00000513061000ef",
        INIT_71 => X"00000013029000ef00100513031000ef00000513039000ef00000513041000ef",
        INIT_72 => X"0201041300812c2300112e23fe01011300008067020101130181240301c12083",
        INIT_73 => X"0ff7f593fe8427830ff7f713fec42783fed42023fec42223feb42423fea42623",
        INIT_74 => X"00050713fe8ff0ef00070513000786930ff7f793fe0427830ff7f613fe442783",
        INIT_75 => X"0ff7f613fe4427830ff7f593fe8427830ff7f713fec427830cf70e6300100793",
        INIT_76 => X"0af70663001007930005071394dff0ef00070513000786930ff7f793fe042783",
        INIT_77 => X"0ff7f793fe0427830ff7f613fe4427830ff7f593fe8427830ff7f713fec42783",
        INIT_78 => X"0ff7f713fec4278306f70e630010079300050713aa5ff0ef0007051300078693",
        INIT_79 => X"00070513000786930ff7f793fe0427830ff7f613fe4427830ff7f593fe842783",
        INIT_7A => X"0ff7f593fe8427830ff7f713fec4278304f706630010079300050713bc9ff0ef",
        INIT_7B => X"0200006fd09ff0ef00070513000786930ff7f793fe0427830ff7f613fe442783",
        INIT_7C => X"01c12083000000130080006f000000130100006f000000130180006f00000013",
        INIT_7D => X"fea426230201041300812c2300112e23fe010113000080670201011301812403",
        INIT_7E => X"00812c2300112e23fe01011300008067020101130181240301c1208300000013",
        INIT_7F => X"820007b7fef424230ff7f7930107d7930007a78300878793820007b702010413",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"fe4425830030061300000693fef422230ff7f7930087d7930007a78300878793",
        INIT_01 => X"0187d713fe042783fea420230c9000ef08c0006ffe042623ca4ff0effe842503",
        INIT_02 => X"fe04278396e7aa23000047b70ff7f7130107d793fe04278396e7a823000047b7",
        INIT_03 => X"96e7ae23000047b70ff7f713fe04278396e7ac23000047b70ff7f7130087d793",
        INIT_04 => X"97c7a783000047b79787a603000047b79747a583000047b79707a703000047b7",
        INIT_05 => X"000017b7fec42703fef4262300178793fec42783da9ff0ef0007051300078693",
        INIT_06 => X"030104130281242302112623fd0101130000006fcedff0eff6e7f6e3ea578793",
        INIT_07 => X"fec4270300078a630017f793fd8427830380006ffe042623fcb42c23fca42e23",
        INIT_08 => X"0017d793fd842783fcf42e2300179793fdc42783fef4262300f707b3fdc42783",
        INIT_09 => X"030101130281240302c1208300078513fec42783fc0794e3fd842783fcf42c23",
        INIT_0A => X"fe042623fcb42c23fca42e23030104130281242302112623fd01011300008067",
        INIT_0B => X"00f717b3fd842703fe842783fef42423fff78793fe842783fef4242301000793",
        INIT_0C => X"fcf42e2340f707b3fdc4270300f717b3fd842703fe84278302f76c63fdc42703",
        INIT_0D => X"fe842783fef4262300e787b3fec427830007871300f717b300100713fe842783",
        INIT_0E => X"fe01011300008067030101130281240302c1208300078513fec42783fa0794e3",
        INIT_0F => X"f49ff0effec42503fe842583feb42423fea426230201041300812c2300112e23",
        INIT_10 => X"fef4262340e787b3fec4278300050713ec5ff0ef00078513fe84258300050793",
        INIT_11 => X"00112e23fe01011300008067020101130181240301c1208300078513fec42783",
        INIT_12 => X"0007a703fe842783fec42223feb42423fea426230201041300912a2300812c23",
        INIT_13 => X"00c7a703fe84278300050493f69fe0ef00070513000785930007a783fe442783",
        INIT_14 => X"fe84278300f484b300050793f49fe0ef00070513000785930047a783fe442783",
        INIT_15 => X"00f4873300050793f25fe0ef00070513000785930087a783fe4427830187a703",
        INIT_16 => X"000705130007859300c7a783fe4427830007a703fe84278300e7a023fec42783",
        INIT_17 => X"00070513000785930107a783fe44278300c7a703fe84278300050493ef9fe0ef",
        INIT_18 => X"000785930147a783fe4427830187a703fe84278300f484b300050793ed9fe0ef",
        INIT_19 => X"0007a703fe84278300e7a623fec4278300f4873300050793eb5fe0ef00070513",
        INIT_1A => X"00c7a703fe84278300050493e89fe0ef00070513000785930187a783fe442783",
        INIT_1B => X"fe84278300f484b300050793e69fe0ef000705130007859301c7a783fe442783",
        INIT_1C => X"00f4873300050793e45fe0ef00070513000785930207a783fe4427830187a703",
        INIT_1D => X"00070513000785930007a783fe4427830047a703fe84278300e7ac23fec42783",
        INIT_1E => X"00070513000785930047a783fe4427830107a703fe84278300050493e19fe0ef",
        INIT_1F => X"000785930087a783fe44278301c7a703fe84278300f484b300050793df9fe0ef",
        INIT_20 => X"0047a703fe84278300e7a223fec4278300f4873300050793dd5fe0ef00070513",
        INIT_21 => X"0107a703fe84278300050493da9fe0ef000705130007859300c7a783fe442783",
        INIT_22 => X"fe84278300f484b300050793d89fe0ef00070513000785930107a783fe442783",
        INIT_23 => X"00f4873300050793d65fe0ef00070513000785930147a783fe44278301c7a703",
        INIT_24 => X"00070513000785930187a783fe4427830047a703fe84278300e7a823fec42783",
        INIT_25 => X"000705130007859301c7a783fe4427830107a703fe84278300050493d39fe0ef",
        INIT_26 => X"000785930207a783fe44278301c7a703fe84278300f484b300050793d19fe0ef",
        INIT_27 => X"0087a703fe84278300e7ae23fec4278300f4873300050793cf5fe0ef00070513",
        INIT_28 => X"0147a703fe84278300050493cc9fe0ef00070513000785930007a783fe442783",
        INIT_29 => X"fe84278300f484b300050793ca9fe0ef00070513000785930047a783fe442783",
        INIT_2A => X"00f4873300050793c85fe0ef00070513000785930087a783fe4427830207a703",
        INIT_2B => X"000705130007859300c7a783fe4427830087a703fe84278300e7a423fec42783",
        INIT_2C => X"00070513000785930107a783fe4427830147a703fe84278300050493c59fe0ef",
        INIT_2D => X"000785930147a783fe4427830207a703fe84278300f484b300050793c39fe0ef",
        INIT_2E => X"0087a703fe84278300e7aa23fec4278300f4873300050793c15fe0ef00070513",
        INIT_2F => X"0147a703fe84278300050493be9fe0ef00070513000785930187a783fe442783",
        INIT_30 => X"fe84278300f484b300050793bc9fe0ef000705130007859301c7a783fe442783",
        INIT_31 => X"00f4873300050793ba5fe0ef00070513000785930207a783fe4427830207a703",
        INIT_32 => X"0000806702010113014124830181240301c120830000001302e7a023fec42783",
        INIT_33 => X"fef44703800007b7fef407a3000507930201041300812c2300112e23fe010113",
        INIT_34 => X"00112e23fe01011300008067020101130181240301c120830000001300e7a023",
        INIT_35 => X"0007c703fee4262300178713fec4278301c0006ffea426230201041300812c23",
        INIT_36 => X"01c120830000001300000013fe0790e30007c783fec4278300e7a023800007b7",
        INIT_37 => X"fca42e23030104130281242302112623fd010113000080670201011301812403",
        INIT_38 => X"ffc78793fe842783fef4242300279793fd84278308078263fd842783fcb42c23",
        INIT_39 => X"00f7f793fe442783fef4222300f757b3fdc42703fec427830500006ffef42623",
        INIT_3A => X"800007b7fef401a30007c78300f707b3fe44278300478713000037b7fef42223",
        INIT_3B => X"000037b7fa07d8e3fec42783fef42623ffc78793fec4278300e7a023fe344703",
        INIT_3C => X"00008067030101130281240302c12083000000130080006ff15ff0ef00078513",
        INIT_3D => X"06079863f9c42783fe042623f8a42e23070104130681242306112623f9010113",
        INIT_3E => X"00a005930b40006fec5ff0ef00078513000037b700e7a02303000713800007b7",
        INIT_3F => X"fe442783f8a42e23951ff0eff9c4250300a00593fea422239f9ff0eff9c42503",
        INIT_40 => X"00e7a023fe44270300f707b300271713fa440793fec42703fef4222300f7f793",
        INIT_41 => X"fff78793fec427830440006ffa0796e3f9c42783fef4262300178793fec42783",
        INIT_42 => X"01870713000037370007a78300f707b300271713fa440793fec42703fef42623",
        INIT_43 => X"fa079ee3fec4278300e7a023feb44703800007b7fef405a30007c78300f707b3",
        INIT_44 => X"fd01011300008067070101130681240306c12083e11ff0ef00078513000037b7",
        INIT_45 => X"fdc42703800007b701c0006ffe042623fca42e23030104130281242302112623",
        INIT_46 => X"fce7dee370f787930065b7b7fec42703fef4262300178793fec4278300e7a023",
        INIT_47 => X"00112e23fe01011300008067030101130281240302c120830000001300000013",
        INIT_48 => X"0007a703820007b7fef426230007a78300478793820007b70201041300812c23",
        INIT_49 => X"00e7a023ffe77713820007b70007a703820007b700e7a02300176713820007b7",
        INIT_4A => X"00112623ff01011300008067020101130181240301c1208300078513fec42783",
        INIT_4B => X"0000001300e7a02300376713810007b70007a703810007b70101041300812423",
        INIT_4C => X"010104130081242300112623ff01011300008067010101130081240300c12083",
        INIT_4D => X"00c120830000001300e7a02300176713810007b70007a703810007b7068000ef",
        INIT_4E => X"02c000ef010104130081242300112623ff010113000080670101011300812403",
        INIT_4F => X"0081240300c120830000001300e7a02300276713810007b70007a703810007b7",
        INIT_50 => X"0007a703810007b7010104130081242300112623ff0101130000806701010113",
        INIT_51 => X"00008067010101130081240300c120830000001300e7a023ffc77713810007b7",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;
