--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"004124230031222300112023340111730000001300000013000000131140006f",
        INIT_01 => X"02c1242302b1222302a1202300912e2300812c2300712a230061282300512623",
        INIT_02 => X"05412423053122230521202303112e2303012c2302f12a2302e1282302d12623",
        INIT_03 => X"07c1242307b1222307a1202305912e2305812c2305712a230561282305512623",
        INIT_04 => X"00812203004121830001208300c010ef3420357307f12a2307e1282307d12623",
        INIT_05 => X"02812603024125830201250301c1248301812403014123830101230300c12283",
        INIT_06 => X"04812a03044129830401290303c1288303812803034127830301270302c12683",
        INIT_07 => X"06812e0306412d8306012d0305c12c8305812c0305412b8305012b0304c12a83",
        INIT_08 => X"000001930000011300000093302000733401117307412f8307012f0306c12e83",
        INIT_09 => X"0000059300000513000004930000041300000393000003130000029300000213",
        INIT_0A => X"0000099300000913000008930000081300000793000007130000069300000613",
        INIT_0B => X"00000d9300000d1300000c9300000c1300000b9300000b1300000a9300000a13",
        INIT_0C => X"0000113700018213eef18193deadc1b700000f9300000f1300000e9300000e13",
        INIT_0D => X"30411073fff001133004507330511073e6810113000001173401107300010113",
        INIT_0E => X"00112023ff4101130540006f6f5000ef001000736fd000effe01011300001137",
        INIT_0F => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_10 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_11 => X"0201041300812c2300112e23fe0101130000006f0000006f0000806700c10113",
        INIT_12 => X"fea426236f9000effec4250300500593fef42623fe078793fec42783fea42623",
        INIT_13 => X"0181240301c1208300078513fec42783fea4262375d000effec4250300900593",
        INIT_14 => X"00068713000507930201041300812c2300112e23fe0101130000806702010113",
        INIT_15 => X"000037b7fef4062300070793fef406a300060793fef4072300058793fef407a3",
        INIT_16 => X"64e78923fed44703000037b764e788a3fee44703000037b764e78823fef44703",
        INIT_17 => X"00008067020101130181240301c120830000001364e789a3fec44703000037b7",
        INIT_18 => X"000037b7fef44703fef407a3000507930201041300812c2300112e23fe010113",
        INIT_19 => X"000037b70007871300f717b30037979340d787b300300793000786936547c783",
        INIT_1A => X"02f71463003007936547c703000037b764e7ac23000037b700f707336587a783",
        INIT_1B => X"6407ac23000037b764078a23000037b700e7a0236587270300003737800007b7",
        INIT_1C => X"0000001364e78a23000037b70ff7f713001787936547c783000037b70200006f",
        INIT_1D => X"030104130281242302112623fd01011300008067020101130181240301c12083",
        INIT_1E => X"fdc42783f29ff0ef00078513fef44783fef407a30187d793fdc42783fca42e23",
        INIT_1F => X"fef407a30087d793fdc42783f11ff0ef00078513fef44783fef407a30107d793",
        INIT_20 => X"ee5ff0ef00078513fef44783fef407a3fdc42783ef9ff0ef00078513fef44783",
        INIT_21 => X"0281242302112623fd01011300008067030101130281240302c1208300000013",
        INIT_22 => X"fef4262300f707b3fec4270301879793fdc42783fe042623fca42e2303010413",
        INIT_23 => X"fdc42783fef4262300f707b3fec4270300f777b300ff07b700879713fdc42783",
        INIT_24 => X"fdc42783fef4262300f707b3fec4270300f777b3f0078793000107b70087d713",
        INIT_25 => X"0281240302c1208300078513fec42783fef4262300f707b3fec427030187d793",
        INIT_26 => X"feb42423fea426230201041300812c2300112e23fe0101130000806703010113",
        INIT_27 => X"06f00513e09ff0ef07100513fef4032300070793fef403a30006871300060793",
        INIT_28 => X"fe842503e99ff0effec42503df1ff0ef06600513df9ff0ef06900513e01ff0ef",
        INIT_29 => X"00000013dc9ff0ef00078513fe644783dd5ff0ef00078513fe744783e91ff0ef",
        INIT_2A => X"0201041300812c2300112e23fe01011300008067020101130181240301c12083",
        INIT_2B => X"00088713000806930007861300070593000685130006031300058e1300050e93",
        INIT_2C => X"fef4062300050793fef406a300030793fef40723000e0793fef407a3000e8793",
        INIT_2D => X"fef4042300070793fef404a300068793fef4052300060793fef405a300058793",
        INIT_2E => X"00f70663fea44783fee447030440006f0000079300f70663feb44783fef44703",
        INIT_2F => X"fec4470301c0006f0000079300f70663fe944783fed447030300006f00000793",
        INIT_30 => X"0181240301c1208300078513001007930080006f0000079300f70663fe844783",
        INIT_31 => X"0006871300050793030104130281242302112623fd0101130000806702010113",
        INIT_32 => X"deadc7b7fcf40e2300070793fcf40ea300060793fcf40f2300058793fcf40fa3",
        INIT_33 => X"c85ff0ef00078513fde44783c91ff0ef00078513fdf44783d4dff0efeef78513",
        INIT_34 => X"000037b76517c303000037b76507c703000037b7c79ff0ef00078513fdd44783",
        INIT_35 => X"00078893fdf44503fde44583fdd44603fdc446836537c783000037b76527c803",
        INIT_36 => X"04e7ea6303f0079365c7c703000037b70607826300050793e8dff0ef00030793",
        INIT_37 => X"fdf44703000037b764e78e23000037b70ff7f7130017879365c7c783000037b7",
        INIT_38 => X"000037b764e78923fdd44703000037b764e788a3fde44703000037b764e78823",
        INIT_39 => X"fc00079302078e6365c7c783000037b704c0006f0010079364e789a3fdc44703",
        INIT_3A => X"fef40723fff787930ff7f79300e787b3fef4470365c7c783000037b7fef407a3",
        INIT_3B => X"02c12083000785130000079364078e23000037b7b99ff0ef00078513fee44783",
        INIT_3C => X"0201041300912a2300812c2300112e23fe010113000080670301011302812403",
        INIT_3D => X"00070793fef406a300060793fef4072300058793fef407a30006871300050793",
        INIT_3E => X"fee447830ff7f49300050793a09ff0ef0030051300078593fef44783fef40623",
        INIT_3F => X"fed447830ff7f49300f487b30ff7f793000507939f1ff0ef0050051300078593",
        INIT_40 => X"fec447830ff7f49300f487b30ff7f793000507939d1ff0ef0070051300078593",
        INIT_41 => X"03f7f7930ff7f79300f487b30ff7f793000507939b1ff0ef00b0051300078593",
        INIT_42 => X"fd0101130000806702010113014124830181240301c12083000785130ff7f793",
        INIT_43 => X"fcf40f2300058793fcf40fa30006871300050793030104130281242302112623",
        INIT_44 => X"fdf44783fde44703fdd44603fdc44683fcf40e2300070793fcf40ea300060793",
        INIT_45 => X"fec4278355078713000037b7fef4262300050793ee5ff0ef0007851300070593",
        INIT_46 => X"00f707b300279793fec4278355078713000037b70007c50300f707b300279793",
        INIT_47 => X"000037b70027c60300f707b300279793fec4278355078713000037b70017c583",
        INIT_48 => X"fde44783fdd44803fdc448830037c68300f707b300279793fec4278355078713",
        INIT_49 => X"fef405a303f7f7930ff7f793fec4278304078c6300050793c2dff0effdf44703",
        INIT_4A => X"fde44703000037b764e78823fdf44703000037b79b9ff0ef00078513feb44783",
        INIT_4B => X"0010079364e789a3fdc44703000037b764e78923fdd44703000037b764e788a3",
        INIT_4C => X"00e78023fdf4470300f707b300279793fec4278355078713000037b70780006f",
        INIT_4D => X"000037b700e780a3fde4470300f707b300279793fec4278355078713000037b7",
        INIT_4E => X"55078713000037b700e78123fdd4470300f707b300279793fec4278355078713",
        INIT_4F => X"02c12083000785130000079300e781a3fdc4470300f707b300279793fec42783",
        INIT_50 => X"00050793030104130281242302112623fd010113000080670301011302812403",
        INIT_51 => X"fcf40e2300070793fcf40ea300060793fcf40f2300058793fcf40fa300068713",
        INIT_52 => X"000037b7fef407a3002787930ff7f79340f707b3fdf447036507c783000037b7",
        INIT_53 => X"6527c783000037b7fef40723002787930ff7f79340f707b3fde447036517c783",
        INIT_54 => X"00e7f66300300793fef44703fef406a3002787930ff7f79340f707b3fdd44703",
        INIT_55 => X"fed447030c00006f0000079300e7f66300300793fee447030d40006f00000793",
        INIT_56 => X"0307f7930ff7f79300479793fef447830ac0006f0000079300e7f66300300793",
        INIT_57 => X"0037f793fed44783fef4072300c7f7930ff7f79300279793fee44783fef407a3",
        INIT_58 => X"0ff7f79300f707b3fee4478300078713fef44783fef4062304000793fef406a3",
        INIT_59 => X"00078513feb44783fef405a300e787b3fec447030ff7f79300e787b3fed44703",
        INIT_5A => X"000037b764e788a3fde44703000037b764e78823fdf44703000037b7fc0ff0ef",
        INIT_5B => X"02c12083000785130010079364e789a3fdc44703000037b764e78923fdd44703",
        INIT_5C => X"00050793030104130281242302112623fd010113000080670301011302812403",
        INIT_5D => X"fcf40e2300070793fcf40ea300060793fcf40f2300058793fcf40fa300068713",
        INIT_5E => X"fef44703fef407a3020787930ff7f79340f707b3fde447036517c783000037b7",
        INIT_5F => X"40f707b3fdf447036507c783000037b71080006f0000079300e7f66303f00793",
        INIT_60 => X"00f00793fee44703fef40723fe8787930ff7f79340e787b3fef447030ff7f793",
        INIT_61 => X"0ff7f79340f707b3fdd447036527c783000037b70cc0006f0000079300e7f663",
        INIT_62 => X"00e7f66300f00793fed44703fef406a3fe8787930ff7f79340e787b3fef44703",
        INIT_63 => X"fec447030ff7f79303f7f793fef44783fef40623f80007930900006f00000793",
        INIT_64 => X"0ff7f71300479793fee44783e70ff0ef00078513fec44783fef4062300e787b3",
        INIT_65 => X"e44ff0ef00078513fec44783fef4062300f707b30ff7f79300f7f793fed44783",
        INIT_66 => X"fdd44703000037b764e788a3fde44703000037b764e78823fdf44703000037b7",
        INIT_67 => X"0281240302c12083000785130010079364e789a3fdc44703000037b764e78923",
        INIT_68 => X"0006871300050793030104130281242302112623fd0101130000806703010113",
        INIT_69 => X"000037b7fcf40e2300070793fcf40ea300060793fcf40f2300058793fcf40fa3",
        INIT_6A => X"fec4278301079713fdf44783fef42623fe0007b706f71a63fdc447036537c783",
        INIT_6B => X"fec42503fef4262300f707b3fdd4478300f7073300879793fde4478300f70733",
        INIT_6C => X"000037b764e788a3fde44703000037b764e78823fdf44703000037b7e30ff0ef",
        INIT_6D => X"000007930080006f0010079364e789a3fdc44703000037b764e78923fdd44703",
        INIT_6E => X"0281242302112623fd01011300008067030101130281240302c1208300078513",
        INIT_6F => X"fcf40ea300060793fcf40f2300058793fcf40fa3000687130005079303010413",
        INIT_70 => X"fdd4478300f7073301079793fde4478301879713fdf44783fcf40e2300070793",
        INIT_71 => X"feb44783fef405a3fff00793fef4262300f707b3fdc4478300f7073300879793",
        INIT_72 => X"030101130281240302c1208300000013d64ff0effec42503cbcff0ef00078513",
        INIT_73 => X"000037b7fef407a3fc0007930201041300812c2300112e23fe01011300008067",
        INIT_74 => X"000037b7c68ff0ef00078513fee44783fef4072300e787b3fef4470365c7c783",
        INIT_75 => X"cf4ff0effe842503fef4242300100793d04ff0effe842503fe04242364078e23",
        INIT_76 => X"0281242302112623fd01011300008067020101130181240301c1208300000013",
        INIT_77 => X"fef407230107d793fdc42783fef407a30187d793fdc42783fca42e2303010413",
        INIT_78 => X"0ff7f7130187d793fdc42783fef40623fdc42783fef406a30087d793fdc42783",
        INIT_79 => X"0ff6f693fdc426830ff7f7930087d793fdc427830ff7f5930107d793fdc42783",
        INIT_7A => X"fdc4278310f70c63001007930007871300050793ee0ff0ef0007051300078613",
        INIT_7B => X"0ff7f7930087d793fdc427830ff7f5930107d793fdc427830ff7f7130187d793",
        INIT_7C => X"0010079300078713000507938cdff0ef00070513000786130ff6f693fdc42683",
        INIT_7D => X"fdc427830ff7f5930107d793fdc427830ff7f7130187d793fdc427830cf70c63",
        INIT_7E => X"00050793a35ff0ef00070513000786130ff6f693fdc426830ff7f7930087d793",
        INIT_7F => X"0107d793fdc427830ff7f7130187d793fdc4278308f70c630010079300078713",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"00070513000786130ff6f693fdc426830ff7f7930087d793fdc427830ff7f593",
        INIT_01 => X"0ff7f7130187d793fdc4278304f70c63001007930007871300050793b6dff0ef",
        INIT_02 => X"0ff6f693fdc426830ff7f7930087d793fdc427830ff7f5930107d793fdc42783",
        INIT_03 => X"0100006f000000130180006f000000130200006fca1ff0ef0007051300078613",
        INIT_04 => X"fe01011300008067030101130281240302c12083000000130080006f00000013",
        INIT_05 => X"020101130181240301c1208300000013fea426230201041300812c2300112e23",
        INIT_06 => X"0007a78300878793820007b70201041300812c2300112e23fe01011300008067",
        INIT_07 => X"fee44783fef406a30087d7930007a78300878793820007b7fef407230107d793",
        INIT_08 => X"0200006ffe0407a3bb4ff0ef00078513000705930030061300000693fed44703",
        INIT_09 => X"fef44703fef407a300178793fef44783da9ff0effe842503fea42423059000ef",
        INIT_0A => X"030104130281242302112623fd0101130000006fd1dff0effce7fee303f00793",
        INIT_0B => X"fec4270300078a630017f793fd8427830380006ffe042623fcb42c23fca42e23",
        INIT_0C => X"0017d793fd842783fcf42e2300179793fdc42783fef4262300f707b3fdc42783",
        INIT_0D => X"030101130281240302c1208300078513fec42783fc0794e3fd842783fcf42c23",
        INIT_0E => X"fe042623fcb42c23fca42e23030104130281242302112623fd01011300008067",
        INIT_0F => X"00f717b3fd842703fe842783fef42423fff78793fe842783fef4242301000793",
        INIT_10 => X"fcf42e2340f707b3fdc4270300f717b3fd842703fe84278302f76c63fdc42703",
        INIT_11 => X"fe842783fef4262300e787b3fec427830007871300f717b300100713fe842783",
        INIT_12 => X"fe01011300008067030101130281240302c1208300078513fec42783fa0794e3",
        INIT_13 => X"f49ff0effec42503fe842583feb42423fea426230201041300812c2300112e23",
        INIT_14 => X"fef4262340e787b3fec4278300050713ec5ff0ef00078513fe84258300050793",
        INIT_15 => X"00112e23fe01011300008067020101130181240301c1208300078513fec42783",
        INIT_16 => X"0007a703fe842783fec42223feb42423fea426230201041300912a2300812c23",
        INIT_17 => X"00c7a703fe84278300050493ee9fe0ef00070513000785930007a783fe442783",
        INIT_18 => X"fe84278300f484b300050793ec9fe0ef00070513000785930047a783fe442783",
        INIT_19 => X"00f4873300050793ea5fe0ef00070513000785930087a783fe4427830187a703",
        INIT_1A => X"000705130007859300c7a783fe4427830007a703fe84278300e7a023fec42783",
        INIT_1B => X"00070513000785930107a783fe44278300c7a703fe84278300050493e79fe0ef",
        INIT_1C => X"000785930147a783fe4427830187a703fe84278300f484b300050793e59fe0ef",
        INIT_1D => X"0007a703fe84278300e7a623fec4278300f4873300050793e35fe0ef00070513",
        INIT_1E => X"00c7a703fe84278300050493e09fe0ef00070513000785930187a783fe442783",
        INIT_1F => X"fe84278300f484b300050793de9fe0ef000705130007859301c7a783fe442783",
        INIT_20 => X"00f4873300050793dc5fe0ef00070513000785930207a783fe4427830187a703",
        INIT_21 => X"00070513000785930007a783fe4427830047a703fe84278300e7ac23fec42783",
        INIT_22 => X"00070513000785930047a783fe4427830107a703fe84278300050493d99fe0ef",
        INIT_23 => X"000785930087a783fe44278301c7a703fe84278300f484b300050793d79fe0ef",
        INIT_24 => X"0047a703fe84278300e7a223fec4278300f4873300050793d55fe0ef00070513",
        INIT_25 => X"0107a703fe84278300050493d29fe0ef000705130007859300c7a783fe442783",
        INIT_26 => X"fe84278300f484b300050793d09fe0ef00070513000785930107a783fe442783",
        INIT_27 => X"00f4873300050793ce5fe0ef00070513000785930147a783fe44278301c7a703",
        INIT_28 => X"00070513000785930187a783fe4427830047a703fe84278300e7a823fec42783",
        INIT_29 => X"000705130007859301c7a783fe4427830107a703fe84278300050493cb9fe0ef",
        INIT_2A => X"000785930207a783fe44278301c7a703fe84278300f484b300050793c99fe0ef",
        INIT_2B => X"0087a703fe84278300e7ae23fec4278300f4873300050793c75fe0ef00070513",
        INIT_2C => X"0147a703fe84278300050493c49fe0ef00070513000785930007a783fe442783",
        INIT_2D => X"fe84278300f484b300050793c29fe0ef00070513000785930047a783fe442783",
        INIT_2E => X"00f4873300050793c05fe0ef00070513000785930087a783fe4427830207a703",
        INIT_2F => X"000705130007859300c7a783fe4427830087a703fe84278300e7a423fec42783",
        INIT_30 => X"00070513000785930107a783fe4427830147a703fe84278300050493bd9fe0ef",
        INIT_31 => X"000785930147a783fe4427830207a703fe84278300f484b300050793bb9fe0ef",
        INIT_32 => X"0087a703fe84278300e7aa23fec4278300f4873300050793b95fe0ef00070513",
        INIT_33 => X"0147a703fe84278300050493b69fe0ef00070513000785930187a783fe442783",
        INIT_34 => X"fe84278300f484b300050793b49fe0ef000705130007859301c7a783fe442783",
        INIT_35 => X"00f4873300050793b25fe0ef00070513000785930207a783fe4427830207a703",
        INIT_36 => X"0000806702010113014124830181240301c120830000001302e7a023fec42783",
        INIT_37 => X"fef44703800007b7fef407a3000507930201041300812c2300112e23fe010113",
        INIT_38 => X"00112e23fe01011300008067020101130181240301c120830000001300e7a023",
        INIT_39 => X"0007c703fee4262300178713fec4278301c0006ffea426230201041300812c23",
        INIT_3A => X"01c120830000001300000013fe0790e30007c783fec4278300e7a023800007b7",
        INIT_3B => X"fca42e23030104130281242302112623fd010113000080670201011301812403",
        INIT_3C => X"ffc78793fe842783fef4242300279793fd84278308078263fd842783fcb42c23",
        INIT_3D => X"00f7f793fe442783fef4222300f757b3fdc42703fec427830500006ffef42623",
        INIT_3E => X"800007b7fef401a30007c78300f707b3fe44278300478713000037b7fef42223",
        INIT_3F => X"000037b7fa07d8e3fec42783fef42623ffc78793fec4278300e7a023fe344703",
        INIT_40 => X"00008067030101130281240302c12083000000130080006ff15ff0ef00078513",
        INIT_41 => X"06079863f9c42783fe042623f8a42e23070104130681242306112623f9010113",
        INIT_42 => X"00a005930b40006fec5ff0ef00078513000037b700e7a02303000713800007b7",
        INIT_43 => X"fe442783f8a42e23951ff0eff9c4250300a00593fea422239f9ff0eff9c42503",
        INIT_44 => X"00e7a023fe44270300f707b300271713fa440793fec42703fef4222300f7f793",
        INIT_45 => X"fff78793fec427830440006ffa0796e3f9c42783fef4262300178793fec42783",
        INIT_46 => X"01870713000037370007a78300f707b300271713fa440793fec42703fef42623",
        INIT_47 => X"fa079ee3fec4278300e7a023feb44703800007b7fef405a30007c78300f707b3",
        INIT_48 => X"fd01011300008067070101130681240306c12083e11ff0ef00078513000037b7",
        INIT_49 => X"fdc42703800007b701c0006ffe042623fca42e23030104130281242302112623",
        INIT_4A => X"fce7dee370f787930065b7b7fec42703fef4262300178793fec4278300e7a023",
        INIT_4B => X"00112e23fe01011300008067030101130281240302c120830000001300000013",
        INIT_4C => X"0007a703820007b7fef426230007a78300478793820007b70201041300812c23",
        INIT_4D => X"00e7a023ffe77713820007b70007a703820007b700e7a02300176713820007b7",
        INIT_4E => X"00112623ff01011300008067020101130181240301c1208300078513fec42783",
        INIT_4F => X"0000001300e7a02300376713810007b70007a703810007b70101041300812423",
        INIT_50 => X"010104130081242300112623ff01011300008067010101130081240300c12083",
        INIT_51 => X"00c120830000001300e7a02300176713810007b70007a703810007b7068000ef",
        INIT_52 => X"02c000ef010104130081242300112623ff010113000080670101011300812403",
        INIT_53 => X"0081240300c120830000001300e7a02300276713810007b70007a703810007b7",
        INIT_54 => X"0007a703810007b7010104130081242300112623ff0101130000806701010113",
        INIT_55 => X"00008067010101130081240300c120830000001300e7a023ffc77713810007b7",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;
