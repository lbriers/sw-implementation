--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     sensor_b - Behavioural
-- Project Name:    sensor_b
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250328   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity sensor_b is
    port(
        clock : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(11 downto 0);
        data_out : out STD_LOGIC_VECTOR(7 downto 0)
    );
end entity sensor_b;

architecture Behavioural of sensor_b is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(11 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(7 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal address_00 : STD_LOGIC_VECTOR(15 downto 0);
    signal data_out_00 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    address_i <= address;
    data_out <= data_out_o;

    address_00 <= "0" & address_i & "000";
    data_out_o <= data_out_00(7 downto 0);
    
    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => x"292e433535412d406e724165644e6f78463035532e2a273938232b2138ff0000",
        INIT_01 => x"0a0c0d0b0f171f1f371e271b1d112b22231e2b1b31391a20262c1e2b203f282e",
        INIT_02 => x"7e6890aaa2514031393027232a2c19301e3c3723240d1d1f322b3f462715080a",
        INIT_03 => x"2f1c161a1f22252b202734313332312c312e342b322a292e3d344c37544f5c5e",
        INIT_04 => x"2c2e34282e242823182212172736122e3b2414060a0a0c0d0e2620251d2f1e23",
        INIT_05 => x"343d45302f3f3523373a2b3d3141373f3a454c51838c91b7beac684d3243302b",
        INIT_06 => x"1c1b302b283c1c1e0a0d0b0a0f151820241e4f2b1a2d2c1b271d212b21214b2b",
        INIT_07 => x"38373e3a3f3c453d48969194ab8f6544472e463e32302c2e2e232d2523352a0c",
        INIT_08 => x"121824241d332a3b232f2122281b202d2828263a46443a482d2f5342303b3a31",
        INIT_09 => x"ab93715d4c4236404b3c32352e2f3e31232c252b15131f201c242f27220d0f0c",
        INIT_0a => x"2c291e232330273130403e30482f2f43362e3d38372b2643455f47594e537599",
        INIT_0b => x"45322d3d2a323e2c33150b1c222725331e1811110e0c0e26221d262e4b3b2c18",
        INIT_0c => x"373d2d343b382d3d3b4333394b3e4e41555a5f6c9c8f6e7969544e4861483c2f",
        INIT_0d => x"1e28232d302b1b0e100f0f191d27242a2e42582b15121e1e233027382f383d45",
        INIT_0e => x"3e4e435742596a97998c7c83797955534c57413840314f253a3d2835282f200e",
        INIT_0f => x"1a292633373b576d462617212e2833343a354342422935302d3a232642424c38",
        INIT_10 => x"76687e625741424e4e4440263636252527303117111e2224322b23200d0e0c0f",
        INIT_11 => x"203432595838383a423d3a453a323225283c433f3d584949614c679bb9958388",
        INIT_12 => x"343629282630442d171a29212d261e2019100f0e12152a2c2b2d48595254382a",
        INIT_13 => x"42413a392a3c4546474f54494259546085a58d817d7b6865585043524d4c283e",
        INIT_14 => x"1d2131281e1b11100e0f1e2b24272b36414e49453235332c4a58443737434049",
        INIT_15 => x"575054596a839c9991a29b7c6454534d57594f43364233202f272c373a172026",
        INIT_16 => x"2e2f2a2e39344a484739343a2a38374e3a36364c6a50473a37303e434f586d5d",
        INIT_17 => x"88886353585a605f55553d42312e29312e43101921252522351c141315141919",
        INIT_18 => x"2d332c3636343e3f42695b503d3a2d3d4e4d666a556b565d618d96978e8d8781",
        INIT_19 => x"404531362e324d181726272a20251b171411131a1f292f32363f39433a39342b",
        INIT_1a => x"4f42435d564c5c646a6167566573898d9aa2857a8b9eaa78535e5760524d524e",
        INIT_1b => x"2a2a31151216151013152b302d3834354743403822342f38334031553649685d",
        INIT_1c => x"5b6672878395ae92859ab3ab7150555f6d6a6a71594942333c362131161a262e",
        INIT_1d => x"24273b3b4460574149395832493d3f3c57366e605c4b454b7e6a4d586b766e81",
        INIT_1e => x"9b735562757d84997f6b53383043372f301d1c283c3920271616111714131a28",
        INIT_1f => x"3b3f4e493c58416660684d4a5b8c775d636e7d6b775e6f6e84a0b0ac9daca99e",
        INIT_20 => x"3e33352438311c1c2b3d3726281513131210161a2b312a303f5a6358464d3f43",
        INIT_21 => x"4e678d7d6763768874816475798ab7c8b8aeb8b09d897658707499a0a37d615f",
        INIT_22 => x"2824161211121415192531312d38615c5a5551504b324a533d4354504f646f48",
        INIT_23 => x"78798ebed2c3b3bbbaaa8f70647894bbaeb1845e4c33291a1a3734171c2c3736",
        INIT_24 => x"323a36504b7272623b3f343f31383343474b5a6852506a8a7a6b618197818669",
        INIT_25 => x"6e68758eaab4ae7a6f563f352e28343a15202f413c2f2418111113181c192c28",
        INIT_26 => x"39333f3f46404c6873515461807262608aa08d876a807792afc7b9b2b2b4aaa2",
        INIT_27 => x"5046353d40151d3249352f281b1213161f161d25312c37323e445e5544332c29",
        INIT_28 => x"5b75685e6489ad8c866d796f9dadb5b1b6b2ae928a726a8a91a9aabd8161735e",
        INIT_29 => x"2b201516191b1621212e3033334137544b542e32273d45342c4f3d4e6c665959",
        INIT_2a => x"69aebcb6b3b9b1a699886c6e7a9db1acae877083675765654f3516202d403b30",
        INIT_2b => x"3a373634455459373834414742334b37726a66575764775d5f5f85a4847d6467",
        INIT_2c => x"6f7897ab9b8c7b6f7c6353565c4a34151e28584835281f171a171d1e261d2f34",
        INIT_2d => x"473f2d5a39706b5d554e647f6a5e567884737d5e6273abb6b1a7b0b1a39e9674",
        INIT_2e => x"6d514540141926503e2d252016131c1d221b202e2b303b2a2540595d3242294c",
        INIT_2f => x"7866555c7c8a7e7e5e6878a4aaa5aeadac997877526d8b8daba297876772746d",
        INIT_30 => x"1e1b101e101b1a2929242f2f1e322a40483a3a3043373333363c4f615a4e435b",
        INIT_31 => x"9ba99ba8b586868f8a5b5694918e8d88746673837569594d390d1926403a2c24",
        INIT_32 => x"31362b2c3f48373b2d3331363c423e464f484b4059625d4a6184928a82567074",
        INIT_33 => x"88898e7d72716075827568555043121b2433342f211e1a191317212126221b32",
        INIT_34 => x"44464c444748404a4053564f485c818d98854c686aaba7a1ae7b8fa88d854c5f",
        INIT_35 => x"63524812181d272f322923181b181a121a1e2c1c2f324433354b573d3b333d42",
        INIT_36 => x"4e465e828e8c876172779a9b97799093a18a7350627b85816d5e6b63707c7e6b",
        INIT_37 => x"1d1a1a1412251d2e232f332c2e45545e413c3c3d423a3a33394d403e3637555a",
        INIT_38 => x"8f7c72908988785e4557716d6a665f4c5655636b5e534d3b14191922312b2136",
        INIT_39 => x"344a4444433340373b45372e3b33475043322e575056475e7b8888775d4e688d",
        INIT_3a => x"535255535d4d3a495549554639161d20293031282a21161816181d1429232e3a",
        INIT_3b => x"2f3c37393b49364a4f524648636b717c57584c556b714f74757c79694741584e",
        INIT_3c => x"503b171d20252c2b18211d13150f141c1c10262524342f333a3028333a393833",
        INIT_3d => x"424e5a667152534743645138534e5a4f363c413a3c554e3a2d4a4a353c2d3637",
        INIT_3e => x"1816110f1c181e3025322627292f342f2d503b3c2b323c344143482e394b4c4b",
        INIT_3f => x"60585757524637283c3c36302b3733272a2a2f3338332f121c1720252e21241e",
        INIT_40 => x"212e39372a342f3b28312b333b474542483640464e48434b453c3e4e4b444244",
        INIT_41 => x"27392d441c1d2c3638412c31101f2c2f2b231b211f171414131c181229302926",
        INIT_42 => x"343b5441525e5b635f49534154434949474b45375b4b5049413f4233393b3629",
        INIT_43 => x"19131d1d1c2a32382d1d0813111e2519171f30242e262a323a333c2e49423739",
        INIT_44 => x"2129342b34464a4d3a2e394240453f37333a535c373424273039342a212f3f31",
        INIT_45 => x"100e16191f171933243642382e3a3b4130282220172a2e322c2e2d3c59714c35",
        INIT_46 => x"4c48443322293e31312a2d2c2936373f30292828241d142a2926232c3e36190c",
        INIT_47 => x"2d5035293629382f38323134494746484e4f71453b423a334c55545954575650",
        INIT_48 => x"201c20191e332a282731280f2335333a40453a25070d0f1219221f242d29381f",
        INIT_49 => x"424937414a4f46755344372c485150535c55564d4e543f4a4a413a2e2c282818",
        INIT_4a => x"0b202726352e2b341d060e100f171b1b2c2b3631404244342e1a183038382b32",
        INIT_4b => x"444544484d524e4c464c4d3b3841453d292428261e2623232d3432322d292726",
        INIT_4c => x"090d181c171929332d373e3a432e1d23371b2c271d2a3a3f484b3b3b686a342f",
        INIT_4d => x"413934383637372c131f1f1c18332e382f373126240e1d262e2e373324160b0e",
        INIT_4e => x"2b29321c392c152931302225252f444c46427636423a29393c41494f50403736",
        INIT_4f => x"1c1d281b392c2b3c2c21191f20292c3031240c090a080a1728181b293e31392d",
        INIT_50 => x"2e2e2920274e3c59403738363131242a3c384040404344313638312f24161424",
        INIT_51 => x"1611161823201e120b0d080b15251d1923351f2e40242929212d181e2219202b",
        INIT_52 => x"39382c2926382c443438423e3e43373f26111117171f1d171d182b2b2c321b10",
        INIT_53 => x"0f18211e1c22380f2b311e1e182a1f171a1b13151a1d242523253b36394c2923",
        INIT_54 => x"3729302e2324141227231a14101b21201a1f271c11110c0a1d1d18150d100804",
        INIT_55 => x"33271c1b2525191c1916141f212b231d192b39382224322f211c1c152018383e",
        INIT_56 => x"2a1b211d261c0b110b1015080514180d13091207050f131c1914273e242c1a28",
        INIT_57 => x"161b19100d1a0b1b2c43251d2e23222c2b2b272c2b2931393737211b08132728",
        INIT_58 => x"0604080b0a18070c090412191f1e1e17222a1e18271c1f2a3427322612122022",
        INIT_59 => x"1c2628252e2726322f2e1e27352f331c271109231a1d1f2a20211c160f120907",
        INIT_5a => x"181c211d1c332c2b2425160b0a2e1823262310121d1b1219181119141017211b",
        INIT_5b => x"181f1b251e160c10141d0b140c161f25111a1504050b0a0d13180f040d05040d",
        INIT_5c => x"0b15241d1a15122012121b1b0f1411130e110d1229351f232e2c24241f1d1720",
        INIT_5d => x"1b0d1c1a0f151114060b0e080605140a050a02050b111e100f17322a27151c17",
        INIT_5e => x"28150f1b101207131708111127202529393a222a1a151c281f241217151c2b16",
        INIT_5f => x"0c17100b050407030409121d180f141915282011121312171817162b2e473415",
        INIT_60 => x"1820222910181b191511211414181d12171113241e0f0b1f1b100f0a050e0e06",
        INIT_61 => x"191c1412150f26281c1b2a2922111f1f1b1a211a1f131509100e0f0f0b161a10",
        INIT_62 => x"13100c1915121b1f101f171b1c10100d0507111b100a07170707040505040a0f",
        INIT_63 => x"142c132e21271e24222f261b15110e171d14091e14131912162a132723171823",
        INIT_64 => x"0d170d0706080c0c091011150e080a050305050c0b22191516180c1b2b161816",
        INIT_65 => x"1e29360a0f1516120c12100e141e1d190e0c1a1e1f17121b130c070b100d0d0c",
        INIT_66 => x"1b050708060306050a0b15240b1a040a181c2022221b1f291a1f261c1e241e21",
        INIT_67 => x"0d2218141b131813211e1e2021070a1a090c0e0a17252610130f070d0b0b1a11",
        INIT_68 => x"1f05141a0f0c10172d2a11131527342f222418090c1c1f1321070a18231b1917",
        INIT_69 => x"1f1a190f0611010d1318171811130f0b080d0e0c120e07070604080912080b17",
        INIT_6a => x"070b0f281d13240d160f1f1a171d06051521160a0e1810101c171112160f1118",
        INIT_6b => x"0f13120d110b130c0e0b070913070f05121b230d12150414190908091523180d",
        INIT_6c => x"14130b0806040e1015161113110c0c0a1116141e0d05100f15010f0613101516",
        INIT_6d => x"0d0f0e101211081613151214121909101a14271f111619191b1f2f290e0e120e",
        INIT_6e => x"0c0a130e18190d0d1216061114100b09101b081309130d15160a0f04090f0d06",
        INIT_6f => x"0f0a170b1e2416190c0f0d1c1a100f1826150816131910080909090b0e051212",
        INIT_70 => x"06060a12090f0d0c0b060c080b0f0b13070f0e0b0f0f11141a1f0b121215130c",
        INIT_71 => x"0d0f06040d1424171c160f040e110a0b03090b07100d0b0f120a0c121b131711",
        INIT_72 => x"0c03080d0e0f0c12100a0d14171403060b0f12190f120c0e10171b13120f1310",
        INIT_73 => x"040d1b100908030b110e09080e0b0a130c050f11160d0d0b08060c090c080605",
        INIT_74 => x"120b0b0f0d1111151912130f150c03111e160a0b0a100d11100a060d100c0e16",
        INIT_75 => x"00000000000000000000000000000000000000000000000000000e0a0e120d0c",

        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 9, -- 0-72
        READ_WIDTH_B => 9, -- 0-36
        WRITE_WIDTH_A => 9, -- 0-36
        WRITE_WIDTH_B => 9, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => data_out_00,
        DOPADOP => open,
        DOBDO => open,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_ONES(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => C_NULL(3 downto 0),
        DIADI => C_NULL,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => C_NULL(15 downto 0),
        CLKBWRCLK => C_NULL(0),
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => C_NULL(7 downto 0),
        DIBDI => C_NULL,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;
