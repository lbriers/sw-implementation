--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     sensor_r - Behavioural
-- Project Name:    sensor_r
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250328   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity sensor_r is
    port(
        clock : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(11 downto 0);
        data_out : out STD_LOGIC_VECTOR(7 downto 0)
    );
end entity sensor_r;

architecture Behavioural of sensor_r is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(11 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(7 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal address_00 : STD_LOGIC_VECTOR(15 downto 0);
    signal data_out_00 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    address_i <= address;
    data_out <= data_out_o;

    address_00 <= "0" & address_i & "000";
    data_out_o <= data_out_00(7 downto 0);
    
    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => x"33456a52466d486cabd8a1bbb397b1b8815a4e714e43344d48304035450000ff",
        INIT_01 => x"0b0d0e1016212c426a4d473e37374f4a45514b1a51617a976026399e9686462d",
        INIT_02 => x"c1a0c0d1c7765d44564c3c2f3944374d304b514448211f396c624d51351c070b",
        INIT_03 => x"603c3a5549536251235567a0c0812b358fa87844313843565742724b919cb4a8",
        INIT_04 => x"353c4e494b34373a3b4e231a48806551472a190b0b0b0d0f142e2c34557a6050",
        INIT_05 => x"9dcd9f32307f9c604c3a3e62605b45694e91a49fbac3c3dbe1d7916a435f4539",
        INIT_06 => x"142b6a73746f301f0a0e0c0b121f242f37549d6b455559445146586947277e5c",
        INIT_07 => x"68715d4f7358949394cbced4e2cebc907647604e39373e43413c443439595f18",
        INIT_08 => x"131b3033304962886663576e5c5045565a432b616691ba9d3535747c604d3a49",
        INIT_09 => x"ebe2cfcda46450585241384043404e463141494c200f213b3f5c65482b0c100d",
        INIT_0a => x"7c606b524f664533525a7e9d9a4133596a6a534153727e87609d6da39a9db3d4",
        INIT_0b => x"524742534a444d494f1f0a1d363e3c4c2f2112100f0f143136343e6297888172",
        INIT_0c => x"bda6423962917d58465e88a4ab679474b1b8adb8eae3d1dfcfa0615d79565649",
        INIT_0d => x"223f3f3d3d3522100e0f1421273c3f436b90a497a59a6f776a504a48386a6b9d",
        INIT_0e => x"98a7729374c0cad8e2e9e6e9d7d394675a786a7c8757714f799264574f5d220d",
        INIT_0f => x"22343b4d517ba2b9b9d0ab635d505c5441407876acc0a84139729481624a6684",
        INIT_10 => x"d6c6d09b7552759abcb07f596e9aa58b6f6b5a1e10243f453b312b28110c0d14",
        INIT_11 => x"515e528b8a50455f699ec3ab493c6895855a4a608ca39d7d9881c1e9f2e4e2ec",
        INIT_12 => x"5e6c95b7967c79482313293d4e3223241b0f0d0f171d34404547769497c3cca1",
        INIT_13 => x"9b5541698f8e624d6da0a19e859b9ab6d0e5eae2d9d9c8b9936f5792a3ba967d",
        INIT_14 => x"303a413322170c0e0f142535394245506e8da7a56c4d5845607f634b5f6a99be",
        INIT_15 => x"9c9093a1b9cfdcebe7f4edd2b99068618b887c7b706d6d84a9865d60621c1624",
        INIT_16 => x"384447474c56728a705547504553626a506a669bae9564416f9a8862577cb4ac",
        INIT_17 => x"dccf9a6c6e787878747d696c65766d6758501716252d29324524151013151e1f",
        INIT_18 => x"685861705d51929ab2c8b374487194836c5a92b9abb18f929bd4e2dde2ebebe2",
        INIT_19 => x"7463586369695e1d152b2e2e21261d19120e141e2532454e4f55605756567372",
        INIT_1a => x"7a5078bc996a6d9ac1baac8c96aad0dae2ede1e1e7e2e5a96e7b798173717487",
        INIT_1b => x"2e272d1311131311171c34454a51607e757c868e71796a79736751b08db7beae",
        INIT_1c => x"949db3d4d2dceee3dfe0e2db9c6f798293908d8ea5936c5e66766c611a182a35",
        INIT_1d => x"3944545a8a93a0977a5470588072605cab86d5b3ae7b567fdbab6b6da8cec3c6",
        INIT_1e => x"c89e7389a2abacb694a786746a7e7473681f192c443d212816140c1515182131",
        INIT_1f => x"455c7161569575b8aeb47d5c88d8b27677acdacfca9babb3d3e1e8ebdee9dec8",
        INIT_20 => x"8a7c81776d5e20192b4537262914100f10111a203342454e597e96a18f6f544f",
        INIT_21 => x"5f8fd0b5847bb3e0d7d5a1b3c1d8ecf0eae1e7dccec7af7f9ba0c7cdcb9a9b9a",
        INIT_22 => x"2522130f0d0f151a202d434b4c4e77808e8b7364563e6375535a8384b0bebd7a",
        INIT_23 => x"b9c2daecf0e8d9e0ddd2c69f7f96aed6cbd2a59193879c93919c721a192b4035",
        INIT_24 => x"4c5a4d65679ba18857554a5d564e476b7ab2b8b5835f90ccb18f82bae5dbd5a6",
        INIT_25 => x"947f91a7bdc6c59a989b89aca4848577171d2e4a3a261e140f0e111920203439",
        INIT_26 => x"5d5a55507571a3b9bb775f89c8ab8c88c0e5dfd2a6c3c0dfe1ead9d2d2d4cbcc",
        INIT_27 => x"98886c646e151a315234231e15111113201b242d4047565361739993745b504f",
        INIT_28 => x"86bc9f8d8fc4f3dcd1aab9afe7e2ddd2d4d2d4bfc3a68bb0b6beb9d49c8bc1a4",
        INIT_29 => x"201812171b1d1b2b2c3d4854576d719a918f625f516c744f41836c9fbbaf7b61",
        INIT_2a => x"a3f3efe0d7d9d4d0ccc39e8c99b9bfb9c9a79bc8a77f8f8e7a621a1c34563f27",
        INIT_2b => x"5c575d6a8091956a605474785d4b7b64c5bbb17b6092b6919189c3f0d6cda5a7",
        INIT_2c => x"8192aabbb4b6ab90a0896d6e78695514203c7a56312016131e1b1f23322d3f4b",
        INIT_2d => x"7155438661bbb19d775a94bc9f907eb2cfc6cea0a3b0efe8ded2dbddd1c9c094",
        INIT_2e => x"7a635d5c15233e75532d1f191418201e2627313f4454594f54758c8d5b624476",
        INIT_2f => x"b29d8881b1cfcbc999a4b9e7dcd5e1e3e3cca09a6b81b0b0ccc8c6b5828a8f7d",
        INIT_30 => x"191c16221220263c3d3f55544b686273715e584b6c604b4c5f5c909b906e528e",
        INIT_31 => x"dcdbd0e0f1c1bcbab37470c9cec4bfb79b8091a08371645f511320345d4b2d1f",
        INIT_32 => x"5f67606673705b5c4c5a5c545c6c5f8182766b548c9b967d86b9d3cfc48ba8b8",
        INIT_33 => x"ced5d3bfb6ac818ea28c7357534d0f1b28453e2f1f1b1b1e1719262e3a373758",
        INIT_34 => x"71737c7c867c6c7562868c927487c0d3d2bf809dabe7e0dce4b0c2dbb8b65c7f",
        INIT_35 => x"756662111b28383e382c24171b1a1f1b252f423a545e5d4f5c757e5e5b57646e",
        INIT_36 => x"8b6f88bfd2c4be94a3b4d9d8cfa6bcbcc7b1a5638fc3c2beb0aca98487959488",
        INIT_37 => x"221d1b1a1a312e4441525a536582848560595f747566655c698677705e5b888c",
        INIT_38 => x"d9b6afcfc2baad94588aae9c9ea8b29a8d8a979685716a5f131b23323e352a3c",
        INIT_39 => x"597c7a6a5e4a58556362483d565974827455568c7c8a6c89b5cfc9b99988a7d8",
        INIT_3a => x"787f92a1ab8f84958a6f71625c141d28363b3c3233291a1a1b2028263f405361",
        INIT_3b => x"345255585e6e5871857a736a8da4b3b4908b7e9ac5c88dbabebdb2a78150867b",
        INIT_3c => x"705b151b263136342027211516141c272c27424a504c3b3f4035304758504032",
        INIT_3d => x"657e969693797f7582bd9e6a958d8f7a605948565f817b78698a89797f696b5f",
        INIT_3e => x"191613162421304c4b5b3c292e383a3141794e3e2d33413f4e535a3f546c6b6b",
        INIT_3f => x"9ba09e988c7b583e62696664727b7a645c5c6667625a56111b1e2c3232262a23",
        INIT_40 => x"2531414a423c4a512b362d3c4d5b5b565748545c666569786e62687c7a758276",
        INIT_41 => x"587d70775557575b6166525f132b4049452e2630291b15181a25202343534f3f",
        INIT_42 => x"404b635163706b76775b665c776d77797a7e7465848990857c7875544f5d5a55",
        INIT_43 => x"4614232b303f434c412b0f15172730242938504b472d323e585b493b62483e43",
        INIT_44 => x"41515e596c8a9496795b6e7872746a604d4f6f735c5958535c5d515350546258",
        INIT_45 => x"141520262c2a34514850525351565868494523211f353b3d343a434f7598674f",
        INIT_46 => x"817c77634945574d494a4b5049535b67564c4a4a4a4614282f332f3e54492511",
        INIT_47 => x"49784d396148563b4b534b4b595659626773a46a636e646183959ca8aaa59185",
        INIT_48 => x"3d3e474040544a474751460f2843474c545b4e310e12151c2631323c4c4b5030",
        INIT_49 => x"8281696e6a7171ab82726557809190949f9e9e928f8f737e7d6f5d4e49434833",
        INIT_4a => x"0c28393d4c4843492d11121215242c2c424a5d5056595d453621274c535a5d75",
        INIT_4b => x"7b827e848c95938f898f947e737373664e47473f343f42434a53515452483d37",
        INIT_4c => x"0b14242b262e455c51535b5856321f334e29373d4c6377859190766c8f9d5c50",
        INIT_4d => x"7e6d605c54534f41232d3137324a46514d574b3a3610283844494f4836241512",
        INIT_4e => x"433a3525583d1625333839586f829a9e8060a95f6a76646c727d898e907f7a78",
        INIT_4f => x"3232392f50443f51433a1b282a384344423117100e0a112335252e445f4c4b3f",
        INIT_50 => x"4a545158749f828b716c74685d5f5c687575838272716e54575a504a3a201d34",
        INIT_51 => x"19121c2835302a1a11110a1121322a293d583d42553c38303c5d221a1a18253a",
        INIT_52 => x"5a635c626f7866b37f626f6f6a67585f3c1a1821273130242a314b4746472e11",
        INIT_53 => x"162332242238583140463e332a563616191b14141a2633394058848a929d5e44",
        INIT_54 => x"65535551453d21172e2f292a212631373337392c12140f0e212b271f12130c09",
        INIT_55 => x"3a3b402223251a1e1b171622273f4e606889a39a5d516b695a525144764f5e69",
        INIT_56 => x"412b2f2b39321d211712180b081723191b0e160b0a161d2d201a3956413d273c",
        INIT_57 => x"151a232d3e545c8a9e97482a443b3d4d4e56434b504f565d5a57382a17253e42",
        INIT_58 => x"09070c13111f0d110d0919222f27232336493120352a374b4d29352a17172323",
        INIT_59 => x"4940424853574c5950504148544f4b2c321a15332d2a2c3b32342f251c1c0c0a",
        INIT_5a => x"212a2c2324474f462e3127161b521f272a2815162221151c292c384a637a7d61",
        INIT_5b => x"353936352a2315171e2c1a231d2831331d251f07080e0e10171d150a12090a14",
        INIT_5c => x"0e2245201e573c231a181e1b111d2126294057769398634543454543413d3842",
        INIT_5d => x"2c1e2c291a1f1b1e09100f12261e2111090e0509111a2f22151d3e484d28231a",
        INIT_5e => x"291515261d1c2268b1b777506d4b3a43524d3a47372a313d2e3425231e263b27",
        INIT_5f => x"193f2d1c0b060a06090f1a312d1319222f4d391811161e2e2527706b38553d19",
        INIT_60 => x"5261595927345137272332242429302722171b332d1d192d281b1a1511141406",
        INIT_61 => x"2d3019191d21403f291e2b2d2d1e2c57492930272b1b180e15131c203b909f60",
        INIT_62 => x"2823222c221b20261c2d2327291b1a170f111b211014252c1209040807091018",
        INIT_63 => x"1b3a1d3631382a312f3c33271e15102e2d2222404152554a554f458851252636",
        INIT_64 => x"172118100e1215160e0f17271e0d09040508091113372d1a1c1e152a40271c1a",
        INIT_65 => x"2d353d0e1c242625262e425f535955574f28272a3932272d2317151417161716",
        INIT_66 => x"280e09060404090a10132737101c0a0f202c3026282530402e273126272e272c",
        INIT_67 => x"415d4d49595746292f33352c2a121c361e18120f1c2a2b1517130c1114141f18",
        INIT_68 => x"2d0e132117111820353318162a424b3c2c30261515242618250d102337353841",
        INIT_69 => x"271e1e1b22280d16181c1b1b1516120e0c1919161b15090806050a0c160e1222",
        INIT_6a => x"070e1c3d3824311e261a261f1b200b091c30291e23312b3247494c51472b2224",
        INIT_6b => x"1216130e120c191314100b0b15081106151f28151f220d182616111626342816",
        INIT_6c => x"19160c0d0807171c21201a1b1d1c25293a3b333d230b12131e12201218141819",
        INIT_6d => x"0f12111214140c1b1b231c1e1e271518252339311b18161b2b3c45391f1c1a14",
        INIT_6e => x"181e26212b362c28292911171c1c110c0f1708140a140e15160a10091216130a",
        INIT_6f => x"191b2513222d2024191a14201c16222c37220d16171c11070c090810170f1d1d",
        INIT_70 => x"171210140b100e0d0c060b060b100c14111b1814161415181e210e17171d2115",
        INIT_71 => x"10100604131e3021211a170a11100a0b040f14111b1b1b1a1d19202a35272821",
        INIT_72 => x"0a04090e0f19161a171012191c19070a11161c2415241d15151e251d15121613",
        INIT_73 => x"0d101a10090a0712181815161614171f1c171d1f28201a110a080e0c0f090604",
        INIT_74 => x"171010141217181d2218241e1c10071d29170c0d0d120e110f0c0d181a111420",
        INIT_75 => x"0000000000000000000000000000000000000000000000000000141416191211",

        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 9, -- 0-72
        READ_WIDTH_B => 9, -- 0-36
        WRITE_WIDTH_A => 9, -- 0-36
        WRITE_WIDTH_B => 9, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
       
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        SBITERR => open,
        DBITERR => open,
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ECCPARITY => open,
        RDADDRECC => open,
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
                
        CLKARDCLK => clock_i,
        ADDRARDADDR => address_00,
        WEA => C_NULL(3 downto 0),
        DIADI => C_NULL,
        DIPADIP => C_NULL(3 downto 0),
        DOADO => data_out_00,
        DOPADOP => open,
        ENARDEN => C_ONES(0),
        REGCEAREGCE => C_NULL(0),
        
        CLKBWRCLK => C_NULL(0),
        ADDRBWRADDR => C_NULL(15 downto 0),
        WEBWE => C_NULL(7 downto 0),
        DIBDI => C_NULL,
        DIPBDIP => C_NULL(3 downto 0),
        DOBDO => open,
        DOPBDOP => open,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0)
    );
                
end Behavioural;
