--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     sensor_g - Behavioural
-- Project Name:    sensor_g
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250328   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity sensor_g is
    port(
        clock : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(11 downto 0);
        data_out : out STD_LOGIC_VECTOR(7 downto 0)
    );
end entity sensor_g;

architecture Behavioural of sensor_g is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(11 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(7 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal address_00 : STD_LOGIC_VECTOR(15 downto 0);
    signal data_out_00 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    address_i <= address;
    data_out <= data_out_o;

    address_00 <= "0" & address_i & "000";
    data_out_o <= data_out_00(7 downto 0);
    
    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => x"2d406a50426b41679cbd88a59e849faa79584c704f4737514b33453b4a00ff00",
        INIT_01 => x"090b0c0c111923416e514c453d3e534d495a50194c5f758f5f2339a08a85472b",
        INIT_02 => x"af8fb0c0b86e5c45554c3e313c493d52355056494c2414366e664c5239210909",
        INIT_03 => x"673e3d5c4e5b6c5722506496b27b283391a3784530333e53513b6f428b8e9c94",
        INIT_04 => x"373f5350513a3c3f41542615457f624f47291c0d09090b0d1028232a55806755",
        INIT_05 => x"91bc972e2e7f9a5f4c3a3a5d5d543b644289968ba8b3b5cdd0c88868445e453a",
        INIT_06 => x"1025666c7973311e090c0a090f171c252b53a16f46565845554d61744c267c5a",
        INIT_07 => x"656e56456f4c868186b7bbc6d3bfad866f415f4d3938424745404a393d5f661b",
        INIT_08 => x"11182829243b5d8a6864576c5b574c5c62462a636886a995323472765e4c3a47",
        INIT_09 => x"d6d0bebf9a5a4b5654483a444944534e37495456220c1e3c405e67492a0a0e0b",
        INIT_0a => x"7a5f6f4f53704d305659718f903a325661634f414f6a757c4d935e9288929dbc",
        INIT_0b => x"544c46544d4752535a21091d3a433e4e301e100f0d0c0f272a272f5a978b806f",
        INIT_0c => x"b19c403a5e85745346587f9aa0528664a1a9a2a5d5d0c1cdbf95565976585c49",
        INIT_0d => x"234445434237210f0e0d101a1c2f3133628da2909f986d7b6850504c356e6690",
        INIT_0e => x"8f9b5c7f61b0b9c8ccd4d3d6c1c1865c5574667a84567653779064565567240d",
        INIT_0f => x"1b282e4041749cafabc3a0595c4f5b57413b786d9eb39e443e6e87795e4b607c",
        INIT_10 => x"bfafbc8c6c4c7290b2a8795d73959d886d7061201025454b43382e2a110c0a10",
        INIT_11 => x"4962568b8e503d5e6191b8a0473f678c7f564a5c879990657f6aacd3decccbd6",
        INIT_12 => x"5f6e8daa8e797b4a27122a42543b2d2a1e0f0d0d131629333737719290b3bd98",
        INIT_13 => x"914c406a8b885e4c689a9995728486a0b9d0d6cdc3c3b3a58466518e96ad8c76",
        INIT_14 => x"36424d3d281a0c0e0d101f2a2b34354c708c9e98674c5f495b816442606792b6",
        INIT_15 => x"9483818da7bcc7d8d3dfd8bda7825b59817d757871706f81a1805d67661f1324",
        INIT_16 => x"2f36363947556f896b5347534955686944676092a38e5d3e6f928260536fa5a0",
        INIT_17 => x"c7bf8c5d64707173737f6c6f65746d6e635819112733343d4d2916101213191a",
        INIT_18 => x"6c5965785e438b8fa4b9a96c446e8a7a675484a8a0a7807b85c0cfc9cad4d5cc",
        INIT_19 => x"72655f6871746820102c3539292c2019120e111a2029363e414c5e555a577276",
        INIT_1a => x"724a71ae8c62658bafaba0797c94bcc7cfd6cdcfd3cdd59a5f6f717a6f707186",
        INIT_1b => x"392f31151113120f13162b3739435a7f74818c93777f707d7a6542a27ba3ada2",
        INIT_1c => x"80839ec1c0c9ddd6d3d0d0cc8e5d6973868685809b8c6e6a6876726c1c132c3c",
        INIT_1d => x"2b334652898b99957d56745f80735a4b9b72c2a4a7724e77cb9c626499bab1b6",
        INIT_1e => x"b98e6279949e9ea57e9d8174697e74766a21142d4a482a2e18140b1513131b29",
        INIT_1f => x"4b5c705b4c8f68a79ca978537ecaa16b6f9bc3bdbc87929cc3d6e1e1d4ded1b9",
        INIT_20 => x"8a7a8580736422142b4d412e2f17100e0f0f161b2c34333e4b77939e8c745854",
        INIT_21 => x"5783c1a37770a0cac6c78c98aac8e0e8e2d8ddd1c2bca3708d96bec4c0879399",
        INIT_22 => x"2d27160f0c0f12161b2735393c4273818e8a75665a4264764f538079a4afb377",
        INIT_23 => x"9aaccae0e6e1d2d9d6c9bd957189a6cec3cb988c9486988d8f9c701c142b4840",
        INIT_24 => x"3a4a43636b9ca08958574e625a4d426872aaadac7f5684bca17e70a6d0ccc68d",
        INIT_25 => x"8a7286a3b9c1c192929b82a59b7e867a18182f51452d22160f0d11171c1b2d2b",
        INIT_26 => x"6561564e776b9aafb471557eba9c7970a9d2d2c38ba0a9cfd5e1d6d0d0d2c5c3",
        INIT_27 => x"968b706a79161631593e2922171111131e161f26333546475c739991745b5355",
        INIT_28 => x"7baf8f7874ace2cebf8f9898d8d8d6d1d3cfd1b8b99c80a7b6bfbad39483bea0",
        INIT_29 => x"221812171a191525242f364148666e958a8f6260556f774d3d836494b1aa7555",
        INIT_2a => x"8de4e5dad5d6cecac2b6927f90b8c2bcc9a190c2a682959581691b173057442a",
        INIT_2b => x"4748586a7c8a956a615673765844795bbbb3ae775286a97f7d70acdfc8ba8a89",
        INIT_2c => x"758aa5bcb7b6a989988972727d6f5c1517327756312016151f191a1d2b233038",
        INIT_2d => x"70513e875bb5ac9c724c89af907f689cbfbbbd87879be0ded9ced5d4c6bcb287",
        INIT_2e => x"7e6864631519336f522e1f1916191e1920202832333f4a4b59778a8c5c644676",
        INIT_2f => x"a590796d9dc2c2b9828ba4d8d2d1dad9d7be918e6078ababcdccc4b67f859283",
        INIT_30 => x"1a1e17210d191f33302d4041436b667472615d506e62494b645b8d9990694584",
        INIT_31 => x"ced0cbd5e5b4ababaa6c6ac6cac5c0b49c7f90a58a766b6759151a2d5b4f3020",
        INIT_32 => x"485a5f6873735f62535f61575f73618282776749828e896f72a6c7c6b87690a5",
        INIT_33 => x"c8cbcab9b5ab7c8ba28d78605a4e101a27494834211c1d1f15151f2631292644",
        INIT_34 => x"797c83828d816d725b7f837f676fa8c7c9b97289a0dad4d0d29fb3cdabb05679",
        INIT_35 => x"7f6e650f192a3c443b2e26181b171b151d2535293f4d534e5e75815f5c5a6c77",
        INIT_36 => x"7e646ea7c6bab7858fa7cccbc196adafbba59d5b89bdbcbaafaeab858999988d",
        INIT_37 => x"241d191515292538303e484b6a888587615a60787869675e6e8c7d735c568485",
        INIT_38 => x"cba6a0c1b5afa28b4d83a49698a2ae9c8f8e9e9b8a7a72611118253644392d3f",
        INIT_39 => x"52807f695e495856635f4439555b78877856538a7886646b9dc6c2b48d7598ca",
        INIT_3a => x"6c718291a38b84988c7177665c121a2939414036372b1b17171b201c32303e50",
        INIT_3b => x"3554555960715a72857777636d8ba9ab897d698ab8ba7da5aaa99f9877427c6d",
        INIT_3c => x"7562121927333a39232a24151410171f231a32363f41383b39312d475a544132",
        INIT_3d => x"5e697d86866a6b5f73aa8957837d806b53503d515e7f756f5a8083747a62655e",
        INIT_3e => x"1a1511121f1d263b354e37282a34362d407d53402f34434251576047576e6d6d",
        INIT_3f => x"8e94938d83755439636d69636f747560555563666159580f1a1f2c3033282c24",
        INIT_40 => x"242f3c4942394a5128332a384857575253434e565e5a5c685d5153625e5c6a62",
        INIT_41 => x"5b8172765557545a68674d58122d434a442e28322a1b151616201b19343f443b",
        INIT_42 => x"353f574455625f67614c5b54736467656161574e7482857a737272514e616059",
        INIT_43 => x"4213242d2f3c424c412a0e1515242b1c1e2a4040442d313b585e47395f40373c",
        INIT_44 => x"40515b51617c82856f4e5e6b676b645d4d5074785f5d5e5a605f525554576254",
        INIT_45 => x"15141d21201d26443f4d54555257596b4948211f1e34393b2f35404d61715b4a",
        INIT_46 => x"75726f5d47465a535052515851565e69564c4a47474212272f312b3b5247210e",
        INIT_47 => x"4c7c4e38664a5a3b4c574e4b5b5b5f6a6e62766163706362839297a1a5a48a78",
        INIT_48 => x"44444e4540524746444d420e2743444751584b2d0b12141a2327272f3e414c32",
        INIT_49 => x"82816a706d756285726e6658829491939d9e9e918e866a76796e6255504d553e",
        INIT_4a => x"0c28383a474641472a0f111014232823353a524d5a5d60473521284c525a6177",
        INIT_4b => x"7b847f848b92928f888e927b7273746c564f514b3d45484a505550514d453e3a",
        INIT_4c => x"0a132429202338524f585f5c57311e344e27363d5066767e8788715e72855251",
        INIT_4d => x"7f70635e575856492d34363d39504a534c564b3c38112a3944464f4835221411",
        INIT_4e => x"463b34255c3f1623333b3c586b7d9598764c87506c76626c717b868c8f7e7a78",
        INIT_4f => x"373940335448445544391c2b2c394347453318100d0810243522253955474c42",
        INIT_50 => x"4f575257729c7c645f7073635c5d5a6573737e817374735a5c5e534f43292438",
        INIT_51 => x"1d131d2838322c1b1110091021342723344f3945583f3a304064241a1918283e",
        INIT_52 => x"5f675e626b77628d6e6673746e6c575537221c252b3736292e37534d4b4b3113",
        INIT_53 => x"121e2e222234532f3f4744372e5f3a191a1a12121a28363b4059868c8e965945",
        INIT_54 => x"675458523e3b281a31332d32292d393e393c3c2f14130e0c202c281f11140d08",
        INIT_55 => x"3b3f47242626191c19161622273f50646c869e955c55716d5b5053435e47606b",
        INIT_56 => x"4b353834433b25281e12170a0716231a1b0d160c091218271e1a35513f3b263f",
        INIT_57 => x"1017243042565c8a9e98462340393b4b4b4f40494d4d535d5b573b301c2a4449",
        INIT_58 => x"08060b13111f0c100e07151c2925231e30472f1e362d3c52522d372a16141f1f",
        INIT_59 => x"463d424a4c514b554a4b3d4352515032371d1938333337473f40392e25240b09",
        INIT_5a => x"1b242b231d424e452c322a191e5924292b2711111d1c111d2b2e394f687f8565",
        INIT_5b => x"323839392f291719212f1f29242f383b242b2606070d0d0f161c1409120a0810",
        INIT_5c => x"0e254c251e3b2d291d171916111d21272f44566d7e8a633f3e3f39383431303d",
        INIT_5d => x"2f212e2c1d221e22070e110f17131c0f0b10060a10182c2416183b4a512a231a",
        INIT_5e => x"261314261e26224b7b89694d69482f3c514f364231232d3e30392b2620283e2a",
        INIT_5f => x"162e24170a0a0e060a101b2e3115161f32533c181117213228234e58415b3f17",
        INIT_60 => x"525c5a5721273c33271d281c2229332c24181d3630201c302a1d1c1713141209",
        INIT_61 => x"2a351b151b2244422a1f2b2e2e1d2541392933292e1c170d1412211c23627e5c",
        INIT_62 => x"251e202c241d20271f3026292b1d1a1710111c2111111a2a120a070a080a1118",
        INIT_63 => x"1d3d1d2f2d322530324238281e150e272c26223b4757514f5b4b2e593f232334",
        INIT_64 => x"1a24190f0d1013180f0e142621110c0606080a121435311c181c152b42291d1b",
        INIT_65 => x"2e363d0d15242b2928354660585557543c1d242b3f36242c2216141318181a19",
        INIT_66 => x"28140f090705090b1114273a121a080e1f2d3228282836473030352225302d34",
        INIT_67 => x"45614b485a594c2d3238392d2a121b2f181612121f2d2e1718140d1212111b14",
        INIT_68 => x"30111320140e16203430181e31494f3c2e31231518252819260c0f2339363742",
        INIT_69 => x"271d1d19161f07141a1e1e1e171814100e13141219150b0b09080b0d170f1324",
        INIT_6a => x"06111f403b2a34161a1528201c200a081c312a1e22322b31474c505649281d21",
        INIT_6b => x"1318181317111a1114110e0c160912061620291622250f1922100a10212d1d0e",
        INIT_6c => x"19160c0c0705171d22211b1b1b1c262b3b3c343c240b11121d07190e1815191b",
        INIT_6d => x"0f11101214140d1b1c261e2021271317252130251216181d2d3f4c3d18111515",
        INIT_6e => x"1b222a25303c322d2e2c12171c1c0c0a121d0b150c16111c1c11160a0b12100a",
        INIT_6f => x"1b1e2a182732231e101516241d1723303a200f1a181d11070c07060e18111f1f",
        INIT_70 => x"19120f140b100f0c0a060d0a0e130f170e0d0d0a0e1012161b210e18181e2416",
        INIT_71 => x"0f0f0706131e3225261d190a0e120a0b020f15131d1d1d1a1d1b232d392a2923",
        INIT_72 => x"0e060c10111f1116120a0d151815030911192027172720161b24271a0f0d1514",
        INIT_73 => x"0e0f1c11090706131a1a1716161418201d191e1f2a221a100a080e0c0c070606",
        INIT_74 => x"130c0c1011181b21241927211c150d1d2411080c0d0f0d11110b0d1b1e161924",
        INIT_75 => x"0000000000000000000000000000000000000000000000000000181113150e0d",

        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 9, -- 0-72
        READ_WIDTH_B => 9, -- 0-36
        WRITE_WIDTH_A => 9, -- 0-36
        WRITE_WIDTH_B => 9, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => data_out_00,
        DOPADOP => open,
        DOBDO => open,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_ONES(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => C_NULL(3 downto 0),
        DIADI => C_NULL,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => C_NULL(15 downto 0),
        CLKBWRCLK => C_NULL(0),
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => C_NULL(7 downto 0),
        DIBDI => C_NULL,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;
